--! @file
--! @brief An almost generic binary to BCD.


----------------------------------------------------------------------------------
-- Engineer (Creator): Jacob Rosén 
-- Engineer (Modifier) : -
--
-- Design Name: binary to BCD coverter
-- Module Name: bin2bcd - Behavioral
-- Project Name: SoundBox
-- Target Devices: Artix 7 
-- 
----------------------------------------------------------------------------------


--! Use of standard library
library IEEE;
--! Use of standard logic arguments
use IEEE.STD_LOGIC_1164.ALL;
--! Use of standard numerical arguments
use IEEE.NUMERIC_STD.ALL;
--! Use of real math arguments to calculate generics.
use IEEE.MATH_REAL.ALL;



entity bin2bcd is
	generic(bits :integer:= 8);
    Port ( bin : in STD_LOGIC_VECTOR (bits-1 downto 0);
           BCD : out STD_LOGIC_VECTOR (bits*2-1 downto 0));
end bin2bcd;

architecture Behavioral of bin2bcd is

component BCD_block
    Port ( in_vector : in STD_LOGIC_VECTOR (3 downto 0);
           out_vector : out STD_LOGIC_VECTOR (3 downto 0));
end component;

constant array_length : integer := bits + integer(floor(real(bits)/real(4)));

type array_type is array (0 to 5 ) of STD_LOGIC_VECTOR(array_length -1 downto 0);
signal temp_vector : array_Type;



begin

generate_loop:
for i in 0 to 4 generate
	gen_temp_values_0: if (i = 0) generate
		temp_vector(0)(array_length -1 downto bits) <= (others => '0');
		temp_vector(0)(bits -1 downto 0) <= bin;
	end generate gen_temp_values_0;


	temp_vector(i+1)(bits-i-4 downto 0) <= temp_vector(i)(bits-i-4 downto 0);

	inst_BCD : BCD_block
		port map (
			in_vector => (temp_vector(i)(bits-i downto bits-i-3)),
			out_vector => (temp_vector(i+1)(bits-i downto bits-i-3))
			);
		
	gen_temp_values : if (i < 3) generate
		temp_vector(i+1)(array_length -1 downto bits+1-i) <= temp_vector(i)(array_length -1 downto bits+1-i);
	
	end generate;
	
	gen_temp_values_4_9 : if i = 3 generate
		inst_BCD : BCD_block
		port map (
				in_vector =>(temp_vector(i)(bits+4-i downto bits+4-i-3)),
				out_vector => (temp_vector(i+1)(bits+4-i downto bits+4-i-3))
				);
	end generate gen_temp_values_4_9;
	
	gen_2nd_row : if i >= 4 generate
		temp_vector(i+1)(array_length -1 downto bits+5-i) <= temp_vector(i)(array_length -1 downto bits+5-i);
		
		
		
		inst_BCD : BCD_block
		port map (
				in_vector =>(temp_vector(i)(bits+4-i downto bits+4-i-3)),
				out_vector => (temp_vector(i+1)(bits+4-i downto bits+4-i-3))
				);
	end generate;
end generate;



BCD(2*bits-1 downto bits+ integer(floor(real(bits)/real(4))) ) <= (others => '0') ;
BCD(bits+ integer(floor(real(bits)/real(4)))-1 downto 0) <= temp_vector(5);



	-- hi : if (i mod 4)  = 0 generate
			-- array_values(i+1) <= array_values(i);
			-- inst_BCD : BCD_block
				-- port map (
					-- in_vector(array_values(i)(bits downto bits-4)),
					-- out_vector(array_values(i+1)(bits downto bits-4))
					-- );	
		-- end generate hi;
		
		-- mid : if (i mod 4)  = 1 generate
			-- array_values(i+1) <= array_values(i);
			-- inst_BCD : BCD_block
				-- port map (
					-- in_vector(array_values(i)(bits -1 downto bits-1-4)),
					-- out_vector(array_values(i+1)(bits -1 downto bits-1-4))
					-- );	
		-- end generate mid;
		
		-- low : if (i mod 4)  = 2 generate
			-- array_values(i+1) <= array_values(i);
			-- inst_BCD : BCD_block
				-- port map (
					-- in_vector(array_values(i)(bits -2 downto bits-2-4)),
					-- out_vector(array_values(i+1)(bits -2 downto bits-2-4))
					-- );	
		-- end generate low;
		
		-- lowhigh : if (i mod 4)  = 3 generate
			-- array_values(i+1) <= array_values(i);
			-- inst_BCD_1 : BCD_block
				-- port map (
					-- in_vector(array_values(i)(bits -3 downto bits-3-4)),
					-- out_vector(array_values(i+1)(bits -3 downto bits-3-4))
					-- );	
			-- inst_BCD_1 : BCD_block
				-- port map (
					-- in_vector(array_values(i)(bits +1 downto bits+1-4)),
					-- out_vector(array_values(i+1)(bits +1 downto bits+1-4))
					-- );	
		-- end generate lowhigh;
		
		-- low : if (i mod 8)  = 4 generate
			-- array_values(i+1) <= array_values(i);
			-- inst_BCD : BCD_block
				-- port map (
					-- in_vector(array_values(i)(bits -2 downto bits-2-4)),
					-- out_vector(array_values(i+1)(bits -2 downto bits-2-4))
					-- );	
		-- end generate low;
		
	
	
	-- if i mod 4 = 0 generate
		

end Behavioral;
